// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.0.240.2
// Netlist written on Mon May  3 15:04:28 2021
//
// Verilog Description of module top_level
//

module top_level (cpu_fpga_bus_a, cpu_fpga_bus_d, cpu_fpga_bus_noe, cpu_fpga_bus_nwe, 
            cpu_fpga_bus_ne1, cpu_fpga_clk, cpu_fpga_int_n, cpu_fpga_rst, 
            fpga_io_gp);   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(5[8:17])
    input [5:0]cpu_fpga_bus_a;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(7[4:18])
    inout [15:0]cpu_fpga_bus_d;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(8[4:18])
    input cpu_fpga_bus_noe;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(9[4:20])
    input cpu_fpga_bus_nwe;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(10[4:20])
    input cpu_fpga_bus_ne1;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(11[4:20])
    input cpu_fpga_clk;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(12[4:16])
    output cpu_fpga_int_n;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(13[4:18])
    input cpu_fpga_rst;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(14[4:16])
    output [7:0]fpga_io_gp;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(15[4:14])
    
    wire cpu_fpga_clk_c /* synthesis is_clock=1, SET_AS_NETWORK=cpu_fpga_clk_c */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(12[4:16])
    
    wire n2907, cpu_fpga_bus_a_c_3, cpu_fpga_bus_a_c_2, cpu_fpga_bus_a_c_1, 
        cpu_fpga_bus_a_c_0, n3119, n3118, n3222, n3117, n3115, n3114, 
        n3113, n3772, n3112, n3111, n3110, n3109, cpu_fpga_bus_nwe_c, 
        cpu_fpga_bus_ne1_c, n2915, cpu_fpga_rst_c, fpga_io_gp_c_7, fpga_io_gp_c_6, 
        fpga_io_gp_c_5, fpga_io_gp_c_4, fpga_io_gp_c_3, fpga_io_gp_c_2, 
        fpga_io_gp_c_1, fpga_io_gp_c_0;
    wire [15:0]\BUFF[15] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[14] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[13] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[12] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[11] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[10] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[9] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[8] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[7] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[6] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[5] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[4] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[3] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[2] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[1] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [15:0]\BUFF[0] ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(26[9:13])
    wire [3:0]address;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(27[9:16])
    
    wire n2661, n3108, n3107, n3106, n3105, n3104, n3103, n3102, 
        VCC_net, n3265, n3085, n3205, n3084, n3083, n3264, n3204, 
        n3082, n3081, n3203, n3080, n3079, n3263, n3202, n3078, 
        n3077, n3201, n3076, n3075, n3262, n3200, n3074, n3073, 
        n3199, n3072, n3070, n3261, n3198, n3069, n3068, n3197, 
        n3067, n3066, n3260, n3196, n3065, n3064, n3195, n3063, 
        n3062, n3259, n3194, n3061, n3060, n3193, n3059, n3058, 
        n3258, n3192, n3057, n3055, n3190, n3054, n3053, n3257, 
        n3189, n3052, n3051, n3188, n3050, n3049, n3256, n3187, 
        n3048, n3047, n3186, n3046, n3045, n3255, n3185, n3044, 
        n3043, n3184, n3042, n3040, n3254, n3183, n3039, n3038, 
        n3182, n3037, n3036, n3253, n3181, n3035, n3034, n3180, 
        n3033, n3032, n3252, n3179, n3031, n3030, n3178, n3029, 
        n3028, n3250, n3177, n3027, n3025, n3175, n3024, n3023, 
        n3249, n3174, n3022, n3021, n3173, n3020, n3019, n3248, 
        n3172, n3018, n3017, n3171, n3016, n3015, n3247, n3170, 
        n3014, n3013, n3169, n3012, n3010, n3246, n3168, n3009, 
        n3008, n3167, n3007, n3006, n3245, n3166, n3005, n3004, 
        n3165, n3003, n3002, n3244, n3164, n3001, n3000, n3163, 
        n2999, n2998, n3243, n3162, n2997, n2995, n3160, n2994, 
        n2993, n3242, n3159, n2992, n2991, n3158, n2990, n2989, 
        n3241, n3157, n2988, n2987, n3156, n2986, n2985, n3240, 
        n3155, n2984, n2983, n3154, n2982, n2980, n3239, n3153, 
        n2979, n2978, n3152, n2977, n2976, n3238, n3151, n2975, 
        n2974, n3150, n2973, n2972, n3237, n3149, n2971, n2970, 
        n3148, n2969, n2968, n3235, n3147, n2967, n2965, n3145, 
        n2964, n2963, n3234, n3144, n2962, n2961, n3143, n2960, 
        n2959, n3233, n3142, n2958, n2957, n3141, n2956, n2955, 
        n3232, n3140, n2954, n2953, n3139, n2952, n2950, n3231, 
        n3138, n2949, n2948, n3137, n2947, n2946, n3230, n3136, 
        n2945, n2944, n3135, n2943, n2942, n3229, n3134, n2941, 
        n2940, n3133, n2939, n2938, n3228, n3132, n2937, n3130, 
        n2934, n3751, n3227, n3129, n2931, n3128, n2930, n3226, 
        n3127, n3126, n2925, n3225, n3125, n2924, n2923, n3124, 
        n2922, n2920, n3224, n3123, n2919, n2918, n3122, n2917, 
        n2916, n3223, n3121, n2914, n2913, n3120, cpu_fpga_bus_d_out_0;
    wire [15:0]cpu_fpga_bus_d_15__N_570;
    
    wire STATE_2__N_297_c_0, cpu_fpga_bus_d_out_1, n3778, n3777, n3776, 
        n3775, n3774, n3773, n3771, n3770, n3769, n3768, n3767, 
        n3766, n3764, n3763, n3762, n3761, n3760, n3759, n3757, 
        n3756, n3755, n3754, n3753, n3752, n3750, n3749, n3748, 
        n3747, n3746, n3745, n3744, n2912, n5, n5_adj_1, n2911, 
        n13, n26, n3765, n2910, n5_adj_2;
    wire [15:0]cpu_fpga_bus_d_15__N_1;
    
    wire GND_net, cpu_fpga_bus_d_15__N_17;
    wire [15:0]fpga_io_gp_7__N_18;
    
    wire n1789, n1790, n1791, n1792, n2655, cpu_fpga_bus_d_out_2, 
        n3758, n2761, cpu_fpga_bus_d_out_3, cpu_fpga_bus_d_out_4, n2760, 
        cpu_fpga_bus_d_out_5, n2909, cpu_fpga_bus_d_out_6, n2692, n2908, 
        cpu_fpga_bus_d_out_7, cpu_fpga_bus_d_out_8, n3534, cpu_fpga_bus_d_out_9, 
        cpu_fpga_clk_c_enable_227, cpu_fpga_clk_c_enable_212, cpu_fpga_bus_d_out_10, 
        cpu_fpga_clk_c_enable_197, cpu_fpga_clk_c_enable_182, cpu_fpga_clk_c_enable_167, 
        cpu_fpga_bus_d_out_11, cpu_fpga_clk_c_enable_152, n2626, cpu_fpga_clk_c_enable_137, 
        cpu_fpga_clk_c_enable_122, cpu_fpga_bus_d_out_12, cpu_fpga_clk_c_enable_107, 
        cpu_fpga_clk_c_enable_92, cpu_fpga_clk_c_enable_77, cpu_fpga_bus_d_out_13, 
        cpu_fpga_clk_c_enable_62, cpu_fpga_clk_c_enable_47, cpu_fpga_clk_c_enable_32, 
        cpu_fpga_bus_d_out_14, cpu_fpga_clk_c_enable_260, n3533, cpu_fpga_clk_c_enable_245, 
        cpu_fpga_bus_d_out_15, cpu_fpga_clk_c_enable_230, n3532;
    
    L6MUX21 i1939 (.D0(n3749), .D1(n3746), .SD(address[2]), .Z(n3750));
    LUT4 i1077_3_lut (.A(\BUFF[10] [5]), .B(\BUFF[11] [5]), .C(address[0]), 
         .Z(n3017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1077_3_lut.init = 16'hcaca;
    BB cpu_fpga_bus_d_pad_9 (.I(cpu_fpga_bus_d_15__N_1[9]), .T(n2626), .B(cpu_fpga_bus_d[9]), 
       .O(cpu_fpga_bus_d_out_9));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    L6MUX21 i1310 (.D0(n3247), .D1(n3248), .SD(\BUFF[0] [2]), .Z(n3250));
    PFUMX i976 (.BLUT(n2909), .ALUT(n2910), .C0(\BUFF[0] [1]), .Z(n2916));
    PFUMX i1937 (.BLUT(n3748), .ALUT(n3747), .C0(address[0]), .Z(n3749));
    BB cpu_fpga_bus_d_pad_10 (.I(cpu_fpga_bus_d_15__N_1[10]), .T(n2626), 
       .B(cpu_fpga_bus_d[10]), .O(cpu_fpga_bus_d_out_10));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    L6MUX21 i1235 (.D0(n3172), .D1(n3173), .SD(address[2]), .Z(n3175));
    BB cpu_fpga_bus_d_pad_11 (.I(cpu_fpga_bus_d_15__N_1[11]), .T(n2626), 
       .B(cpu_fpga_bus_d[11]), .O(cpu_fpga_bus_d_out_11));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    L6MUX21 i1084 (.D0(n3020), .D1(n3021), .SD(address[2]), .Z(n3024));
    L6MUX21 i1085 (.D0(n3022), .D1(n3023), .SD(address[2]), .Z(n3025));
    LUT4 i1076_3_lut (.A(\BUFF[8] [5]), .B(\BUFF[9] [5]), .C(address[0]), 
         .Z(n3016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1076_3_lut.init = 16'hcaca;
    LUT4 i1075_3_lut (.A(\BUFF[6] [5]), .B(\BUFF[7] [5]), .C(address[0]), 
         .Z(n3015)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1075_3_lut.init = 16'hcaca;
    OB cpu_fpga_int_n_pad (.I(GND_net), .O(cpu_fpga_int_n));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(13[4:18])
    BB cpu_fpga_bus_d_pad_12 (.I(cpu_fpga_bus_d_15__N_1[12]), .T(n2626), 
       .B(cpu_fpga_bus_d[12]), .O(cpu_fpga_bus_d_out_12));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    L6MUX21 i1249 (.D0(n3185), .D1(n3186), .SD(address[2]), .Z(n3189));
    L6MUX21 i1250 (.D0(n3187), .D1(n3188), .SD(address[2]), .Z(n3190));
    BB cpu_fpga_bus_d_pad_13 (.I(cpu_fpga_bus_d_15__N_1[13]), .T(n2626), 
       .B(cpu_fpga_bus_d[13]), .O(cpu_fpga_bus_d_out_13));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    L6MUX21 i1099 (.D0(n3035), .D1(n3036), .SD(address[2]), .Z(n3039));
    BB cpu_fpga_bus_d_pad_0 (.I(cpu_fpga_bus_d_15__N_1[0]), .T(n2626), .B(cpu_fpga_bus_d[0]), 
       .O(cpu_fpga_bus_d_out_0));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    L6MUX21 i1100 (.D0(n3037), .D1(n3038), .SD(address[2]), .Z(n3040));
    L6MUX21 i1114 (.D0(n3050), .D1(n3051), .SD(address[2]), .Z(n3054));
    BB cpu_fpga_bus_d_pad_1 (.I(cpu_fpga_bus_d_15__N_1[1]), .T(n2626), .B(cpu_fpga_bus_d[1]), 
       .O(cpu_fpga_bus_d_out_1));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    L6MUX21 i1115 (.D0(n3052), .D1(n3053), .SD(address[2]), .Z(n3055));
    LUT4 i1074_3_lut (.A(\BUFF[4] [5]), .B(\BUFF[5] [5]), .C(address[0]), 
         .Z(n3014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1074_3_lut.init = 16'hcaca;
    BB cpu_fpga_bus_d_pad_14 (.I(cpu_fpga_bus_d_15__N_1[14]), .T(n2626), 
       .B(cpu_fpga_bus_d[14]), .O(cpu_fpga_bus_d_out_14));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    BB cpu_fpga_bus_d_pad_2 (.I(cpu_fpga_bus_d_15__N_1[2]), .T(n2626), .B(cpu_fpga_bus_d[2]), 
       .O(cpu_fpga_bus_d_out_2));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    L6MUX21 i1324 (.D0(n3260), .D1(n3261), .SD(\BUFF[0] [2]), .Z(n3264));
    LUT4 i1073_3_lut (.A(\BUFF[2] [5]), .B(\BUFF[3] [5]), .C(address[0]), 
         .Z(n3013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1073_3_lut.init = 16'hcaca;
    L6MUX21 i1264 (.D0(n3200), .D1(n3201), .SD(address[2]), .Z(n3204));
    LUT4 i1072_3_lut (.A(\BUFF[0] [5]), .B(\BUFF[1] [5]), .C(address[0]), 
         .Z(n3012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1072_3_lut.init = 16'hcaca;
    LUT4 i1177_3_lut (.A(\BUFF[0] [6]), .B(\BUFF[1] [6]), .C(\BUFF[0] [0]), 
         .Z(n3117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1177_3_lut.init = 16'hcaca;
    BB cpu_fpga_bus_d_pad_3 (.I(cpu_fpga_bus_d_15__N_1[3]), .T(n2626), .B(cpu_fpga_bus_d[3]), 
       .O(cpu_fpga_bus_d_out_3));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    PFUMX i1172 (.BLUT(n3106), .ALUT(n3107), .C0(\BUFF[0] [1]), .Z(n3112));
    IB cpu_fpga_rst_pad (.I(cpu_fpga_rst), .O(cpu_fpga_rst_c));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(14[4:16])
    L6MUX21 i1325 (.D0(n3262), .D1(n3263), .SD(\BUFF[0] [2]), .Z(n3265));
    LUT4 i1064_3_lut (.A(\BUFF[14] [6]), .B(\BUFF[15] [6]), .C(address[0]), 
         .Z(n3004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1064_3_lut.init = 16'hcaca;
    FD1P3AX BUFF_12__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i0.GSR = "ENABLED";
    FD1P3AX address_i0_i0 (.D(cpu_fpga_bus_a_c_0), .SP(cpu_fpga_clk_c_enable_230), 
            .CK(cpu_fpga_clk_c), .Q(address[0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam address_i0_i0.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i0.GSR = "ENABLED";
    LUT4 i1063_3_lut (.A(\BUFF[12] [6]), .B(\BUFF[13] [6]), .C(address[0]), 
         .Z(n3003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1063_3_lut.init = 16'hcaca;
    LUT4 i1229_3_lut (.A(\BUFF[14] [15]), .B(\BUFF[15] [15]), .C(address[0]), 
         .Z(n3169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1229_3_lut.init = 16'hcaca;
    PFUMX i1934 (.BLUT(n3745), .ALUT(n3744), .C0(address[0]), .Z(n3746));
    MUX21 i1521 (.D0(n3174), .D1(n3175), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[15]));
    LUT4 i1228_3_lut (.A(\BUFF[12] [15]), .B(\BUFF[13] [15]), .C(address[0]), 
         .Z(n3168)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1228_3_lut.init = 16'hcaca;
    BB cpu_fpga_bus_d_pad_4 (.I(cpu_fpga_bus_d_15__N_1[4]), .T(n2626), .B(cpu_fpga_bus_d[4]), 
       .O(cpu_fpga_bus_d_out_4));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    LUT4 i974_3_lut (.A(\BUFF[14] [2]), .B(\BUFF[15] [2]), .C(\BUFF[0] [0]), 
         .Z(n2914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i974_3_lut.init = 16'hcaca;
    L6MUX21 i1265 (.D0(n3202), .D1(n3203), .SD(address[2]), .Z(n3205));
    PFUMX i1098 (.BLUT(n3033), .ALUT(n3034), .C0(address[1]), .Z(n3038));
    L6MUX21 i979 (.D0(n2915), .D1(n2916), .SD(\BUFF[0] [2]), .Z(n2919));
    L6MUX21 i980 (.D0(n2917), .D1(n2918), .SD(\BUFF[0] [2]), .Z(n2920));
    L6MUX21 i1189 (.D0(n3125), .D1(n3126), .SD(\BUFF[0] [2]), .Z(n3129));
    L6MUX21 i1190 (.D0(n3127), .D1(n3128), .SD(\BUFF[0] [2]), .Z(n3130));
    L6MUX21 i1009 (.D0(n2945), .D1(n2946), .SD(address[2]), .Z(n2949));
    L6MUX21 i1010 (.D0(n2947), .D1(n2948), .SD(address[2]), .Z(n2950));
    L6MUX21 i1294 (.D0(n3230), .D1(n3231), .SD(\BUFF[0] [2]), .Z(n3234));
    L6MUX21 i1204 (.D0(n3140), .D1(n3141), .SD(\BUFF[0] [2]), .Z(n3144));
    L6MUX21 i1295 (.D0(n3232), .D1(n3233), .SD(\BUFF[0] [2]), .Z(n3235));
    L6MUX21 i1205 (.D0(n3142), .D1(n3143), .SD(\BUFF[0] [2]), .Z(n3145));
    LUT4 i1062_3_lut (.A(\BUFF[10] [6]), .B(\BUFF[11] [6]), .C(address[0]), 
         .Z(n3002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1062_3_lut.init = 16'hcaca;
    L6MUX21 i1024 (.D0(n2960), .D1(n2961), .SD(address[2]), .Z(n2964));
    BB cpu_fpga_bus_d_pad_15 (.I(cpu_fpga_bus_d_15__N_1[15]), .T(n2626), 
       .B(cpu_fpga_bus_d[15]), .O(cpu_fpga_bus_d_out_15));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    LUT4 i1061_3_lut (.A(\BUFF[8] [6]), .B(\BUFF[9] [6]), .C(address[0]), 
         .Z(n3001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1061_3_lut.init = 16'hcaca;
    BB cpu_fpga_bus_d_pad_5 (.I(cpu_fpga_bus_d_15__N_1[5]), .T(n2626), .B(cpu_fpga_bus_d[5]), 
       .O(cpu_fpga_bus_d_out_5));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    LUT4 i1060_3_lut (.A(\BUFF[6] [6]), .B(\BUFF[7] [6]), .C(address[0]), 
         .Z(n3000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1060_3_lut.init = 16'hcaca;
    LUT4 i973_3_lut (.A(\BUFF[12] [2]), .B(\BUFF[13] [2]), .C(\BUFF[0] [0]), 
         .Z(n2913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i973_3_lut.init = 16'hcaca;
    LUT4 i1059_3_lut (.A(\BUFF[4] [6]), .B(\BUFF[5] [6]), .C(address[0]), 
         .Z(n2999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1059_3_lut.init = 16'hcaca;
    PFUMX i1173 (.BLUT(n3108), .ALUT(n3109), .C0(\BUFF[0] [1]), .Z(n3113));
    LUT4 i1227_3_lut (.A(\BUFF[10] [15]), .B(\BUFF[11] [15]), .C(address[0]), 
         .Z(n3167)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1227_3_lut.init = 16'hcaca;
    LUT4 i1226_3_lut (.A(\BUFF[8] [15]), .B(\BUFF[9] [15]), .C(address[0]), 
         .Z(n3166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1226_3_lut.init = 16'hcaca;
    LUT4 i1058_3_lut (.A(\BUFF[2] [6]), .B(\BUFF[3] [6]), .C(address[0]), 
         .Z(n2998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1058_3_lut.init = 16'hcaca;
    LUT4 i1057_3_lut (.A(\BUFF[0] [6]), .B(\BUFF[1] [6]), .C(address[0]), 
         .Z(n2997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1057_3_lut.init = 16'hcaca;
    LUT4 i1225_3_lut (.A(\BUFF[6] [15]), .B(\BUFF[7] [15]), .C(address[0]), 
         .Z(n3165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1225_3_lut.init = 16'hcaca;
    LUT4 i1224_3_lut (.A(\BUFF[4] [15]), .B(\BUFF[5] [15]), .C(address[0]), 
         .Z(n3164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1224_3_lut.init = 16'hcaca;
    LUT4 i1304_3_lut (.A(\BUFF[14] [4]), .B(\BUFF[15] [4]), .C(\BUFF[0] [0]), 
         .Z(n3244)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1304_3_lut.init = 16'hcaca;
    BB cpu_fpga_bus_d_pad_6 (.I(cpu_fpga_bus_d_15__N_1[6]), .T(n2626), .B(cpu_fpga_bus_d[6]), 
       .O(cpu_fpga_bus_d_out_6));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    L6MUX21 i1129 (.D0(n3065), .D1(n3066), .SD(address[2]), .Z(n3069));
    LUT4 i972_3_lut (.A(\BUFF[10] [2]), .B(\BUFF[11] [2]), .C(\BUFF[0] [0]), 
         .Z(n2912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i972_3_lut.init = 16'hcaca;
    BB cpu_fpga_bus_d_pad_7 (.I(cpu_fpga_bus_d_15__N_1[7]), .T(n2626), .B(cpu_fpga_bus_d[7]), 
       .O(cpu_fpga_bus_d_out_7));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    LUT4 i1303_3_lut (.A(\BUFF[12] [4]), .B(\BUFF[13] [4]), .C(\BUFF[0] [0]), 
         .Z(n3243)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1303_3_lut.init = 16'hcaca;
    IB cpu_fpga_clk_pad (.I(cpu_fpga_clk), .O(cpu_fpga_clk_c));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(12[4:16])
    LUT4 i971_3_lut (.A(\BUFF[8] [2]), .B(\BUFF[9] [2]), .C(\BUFF[0] [0]), 
         .Z(n2911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i971_3_lut.init = 16'hcaca;
    L6MUX21 i1130 (.D0(n3067), .D1(n3068), .SD(address[2]), .Z(n3070));
    LUT4 i1223_3_lut (.A(\BUFF[2] [15]), .B(\BUFF[3] [15]), .C(address[0]), 
         .Z(n3163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1223_3_lut.init = 16'hcaca;
    L6MUX21 i994 (.D0(n2930), .D1(n2931), .SD(address[2]), .Z(n2934));
    IB cpu_fpga_bus_ne1_pad (.I(cpu_fpga_bus_ne1), .O(cpu_fpga_bus_ne1_c));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(11[4:20])
    L6MUX21 i1144 (.D0(n3080), .D1(n3081), .SD(address[2]), .Z(n3084));
    LUT4 i1222_3_lut (.A(\BUFF[0] [15]), .B(\BUFF[1] [15]), .C(address[0]), 
         .Z(n3162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1222_3_lut.init = 16'hcaca;
    IB cpu_fpga_bus_nwe_pad (.I(cpu_fpga_bus_nwe), .O(cpu_fpga_bus_nwe_c));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(10[4:20])
    IB STATE_2__N_297_pad_0 (.I(cpu_fpga_bus_noe), .O(STATE_2__N_297_c_0));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(9[4:20])
    L6MUX21 i1145 (.D0(n3082), .D1(n3083), .SD(address[2]), .Z(n3085));
    IB cpu_fpga_bus_a_pad_0 (.I(cpu_fpga_bus_a[0]), .O(cpu_fpga_bus_a_c_0));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(7[4:18])
    BB cpu_fpga_bus_d_pad_8 (.I(cpu_fpga_bus_d_15__N_1[8]), .T(n2626), .B(cpu_fpga_bus_d[8]), 
       .O(cpu_fpga_bus_d_out_8));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    LUT4 i970_3_lut (.A(\BUFF[6] [2]), .B(\BUFF[7] [2]), .C(\BUFF[0] [0]), 
         .Z(n2910)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i970_3_lut.init = 16'hcaca;
    IB cpu_fpga_bus_a_pad_1 (.I(cpu_fpga_bus_a[1]), .O(cpu_fpga_bus_a_c_1));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(7[4:18])
    LUT4 i1302_3_lut (.A(\BUFF[10] [4]), .B(\BUFF[11] [4]), .C(\BUFF[0] [0]), 
         .Z(n3242)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1302_3_lut.init = 16'hcaca;
    L6MUX21 i1025 (.D0(n2962), .D1(n2963), .SD(address[2]), .Z(n2965));
    LUT4 i1301_3_lut (.A(\BUFF[8] [4]), .B(\BUFF[9] [4]), .C(\BUFF[0] [0]), 
         .Z(n3241)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1301_3_lut.init = 16'hcaca;
    L6MUX21 i1176 (.D0(n3114), .D1(n3115), .SD(\BUFF[0] [3]), .Z(fpga_io_gp_7__N_18[0]));
    LUT4 i1300_3_lut (.A(\BUFF[6] [4]), .B(\BUFF[7] [4]), .C(\BUFF[0] [0]), 
         .Z(n3240)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1300_3_lut.init = 16'hcaca;
    LUT4 i1299_3_lut (.A(\BUFF[4] [4]), .B(\BUFF[5] [4]), .C(\BUFF[0] [0]), 
         .Z(n3239)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1299_3_lut.init = 16'hcaca;
    LUT4 i1049_3_lut (.A(\BUFF[14] [7]), .B(\BUFF[15] [7]), .C(address[0]), 
         .Z(n2989)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1049_3_lut.init = 16'hcaca;
    L6MUX21 i1039 (.D0(n2975), .D1(n2976), .SD(address[2]), .Z(n2979));
    L6MUX21 i1069 (.D0(n3005), .D1(n3006), .SD(address[2]), .Z(n3009));
    PFUMX i1320 (.BLUT(n3252), .ALUT(n3253), .C0(\BUFF[0] [1]), .Z(n3260));
    LUT4 i1048_3_lut (.A(\BUFF[12] [7]), .B(\BUFF[13] [7]), .C(address[0]), 
         .Z(n2988)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1048_3_lut.init = 16'hcaca;
    L6MUX21 i1040 (.D0(n2977), .D1(n2978), .SD(address[2]), .Z(n2980));
    L6MUX21 i1219 (.D0(n3155), .D1(n3156), .SD(\BUFF[0] [2]), .Z(n3159));
    LUT4 i969_3_lut (.A(\BUFF[4] [2]), .B(\BUFF[5] [2]), .C(\BUFF[0] [0]), 
         .Z(n2909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i969_3_lut.init = 16'hcaca;
    LUT4 i1298_3_lut (.A(\BUFF[2] [4]), .B(\BUFF[3] [4]), .C(\BUFF[0] [0]), 
         .Z(n3238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1298_3_lut.init = 16'hcaca;
    LUT4 i1297_3_lut (.A(\BUFF[0] [4]), .B(\BUFF[1] [4]), .C(\BUFF[0] [0]), 
         .Z(n3237)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1297_3_lut.init = 16'hcaca;
    L6MUX21 i1070 (.D0(n3007), .D1(n3008), .SD(address[2]), .Z(n3010));
    L6MUX21 i1234 (.D0(n3170), .D1(n3171), .SD(address[2]), .Z(n3174));
    L6MUX21 i1220 (.D0(n3157), .D1(n3158), .SD(\BUFF[0] [2]), .Z(n3160));
    LUT4 i1047_3_lut (.A(\BUFF[10] [7]), .B(\BUFF[11] [7]), .C(address[0]), 
         .Z(n2987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1047_3_lut.init = 16'hcaca;
    LUT4 i1046_3_lut (.A(\BUFF[8] [7]), .B(\BUFF[9] [7]), .C(address[0]), 
         .Z(n2986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1046_3_lut.init = 16'hcaca;
    L6MUX21 i1054 (.D0(n2990), .D1(n2991), .SD(address[2]), .Z(n2994));
    LUT4 i1045_3_lut (.A(\BUFF[6] [7]), .B(\BUFF[7] [7]), .C(address[0]), 
         .Z(n2985)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1045_3_lut.init = 16'hcaca;
    LUT4 i1312_3_lut (.A(\BUFF[0] [3]), .B(\BUFF[1] [3]), .C(\BUFF[0] [0]), 
         .Z(n3252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1312_3_lut.init = 16'hcaca;
    L6MUX21 i1309 (.D0(n3245), .D1(n3246), .SD(\BUFF[0] [2]), .Z(n3249));
    L6MUX21 i1055 (.D0(n2992), .D1(n2993), .SD(address[2]), .Z(n2995));
    LUT4 i1044_3_lut (.A(\BUFF[4] [7]), .B(\BUFF[5] [7]), .C(address[0]), 
         .Z(n2984)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1044_3_lut.init = 16'hcaca;
    GSR GSR_INST (.GSR(n2760));
    IB cpu_fpga_bus_a_pad_2 (.I(cpu_fpga_bus_a[2]), .O(cpu_fpga_bus_a_c_2));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(7[4:18])
    IB cpu_fpga_bus_a_pad_3 (.I(cpu_fpga_bus_a[3]), .O(cpu_fpga_bus_a_c_3));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(7[4:18])
    LUT4 i1043_3_lut (.A(\BUFF[2] [7]), .B(\BUFF[3] [7]), .C(address[0]), 
         .Z(n2983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1043_3_lut.init = 16'hcaca;
    LUT4 i1042_3_lut (.A(\BUFF[0] [7]), .B(\BUFF[1] [7]), .C(address[0]), 
         .Z(n2982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1042_3_lut.init = 16'hcaca;
    OB fpga_io_gp_pad_0 (.I(fpga_io_gp_c_0), .O(fpga_io_gp[0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(15[4:14])
    OB fpga_io_gp_pad_1 (.I(fpga_io_gp_c_1), .O(fpga_io_gp[1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(15[4:14])
    PFUMX i977 (.BLUT(n2911), .ALUT(n2912), .C0(\BUFF[0] [1]), .Z(n2917));
    LUT4 i1214_3_lut (.A(\BUFF[14] [1]), .B(\BUFF[15] [1]), .C(\BUFF[0] [0]), 
         .Z(n3154)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1214_3_lut.init = 16'hcaca;
    L6MUX21 i1174 (.D0(n3110), .D1(n3111), .SD(\BUFF[0] [2]), .Z(n3114));
    FD1P3AX BUFF_13__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i0.GSR = "ENABLED";
    OB fpga_io_gp_pad_2 (.I(fpga_io_gp_c_2), .O(fpga_io_gp[2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(15[4:14])
    OB fpga_io_gp_pad_3 (.I(fpga_io_gp_c_3), .O(fpga_io_gp[3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(15[4:14])
    OB fpga_io_gp_pad_4 (.I(fpga_io_gp_c_4), .O(fpga_io_gp[4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(15[4:14])
    LUT4 i1213_3_lut (.A(\BUFF[12] [1]), .B(\BUFF[13] [1]), .C(\BUFF[0] [0]), 
         .Z(n3153)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1213_3_lut.init = 16'hcaca;
    L6MUX21 i1175 (.D0(n3112), .D1(n3113), .SD(\BUFF[0] [2]), .Z(n3115));
    PFUMX i978 (.BLUT(n2913), .ALUT(n2914), .C0(\BUFF[0] [1]), .Z(n2918));
    PFUMX i1185 (.BLUT(n3117), .ALUT(n3118), .C0(\BUFF[0] [1]), .Z(n3125));
    FD1S3IX cpu_fpga_bus_d__i0 (.D(cpu_fpga_bus_d_15__N_570[0]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i0.GSR = "ENABLED";
    OB fpga_io_gp_pad_5 (.I(fpga_io_gp_c_5), .O(fpga_io_gp[5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(15[4:14])
    FD1P3AX BUFF_14__i0_i0 (.D(cpu_fpga_bus_d_out_0), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [0]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i0.GSR = "ENABLED";
    PFUMX i975 (.BLUT(n2907), .ALUT(n2908), .C0(\BUFF[0] [1]), .Z(n2915));
    PFUMX i1186 (.BLUT(n3119), .ALUT(n3120), .C0(\BUFF[0] [1]), .Z(n3126));
    OB fpga_io_gp_pad_6 (.I(fpga_io_gp_c_6), .O(fpga_io_gp[6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(15[4:14])
    OB fpga_io_gp_pad_7 (.I(fpga_io_gp_c_7), .O(fpga_io_gp[7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(15[4:14])
    FD1S3IX i103_278 (.D(n3533), .CK(cpu_fpga_clk_c), .CD(n2761), .Q(cpu_fpga_bus_d_15__N_17));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam i103_278.GSR = "ENABLED";
    PFUMX i1187 (.BLUT(n3121), .ALUT(n3122), .C0(\BUFF[0] [1]), .Z(n3127));
    PFUMX i1188 (.BLUT(n3123), .ALUT(n3124), .C0(\BUFF[0] [1]), .Z(n3128));
    LUT4 i1212_3_lut (.A(\BUFF[10] [1]), .B(\BUFF[11] [1]), .C(\BUFF[0] [0]), 
         .Z(n3152)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1212_3_lut.init = 16'hcaca;
    FD1P3AX BUFF_13__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i1.GSR = "ENABLED";
    LUT4 i1211_3_lut (.A(\BUFF[8] [1]), .B(\BUFF[9] [1]), .C(\BUFF[0] [0]), 
         .Z(n3151)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1211_3_lut.init = 16'hcaca;
    LUT4 i1034_3_lut (.A(\BUFF[14] [8]), .B(\BUFF[15] [8]), .C(address[0]), 
         .Z(n2974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1034_3_lut.init = 16'hcaca;
    FD1P3AX BUFF_13__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_13__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_32), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[13] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_13__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_12__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_47), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[12] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_12__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_11__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_62), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[11] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_11__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_10__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_77), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[10] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_10__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_9__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_92), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[9] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_9__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_8__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_107), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[8] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_8__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_7__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_122), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[7] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_7__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_6__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_137), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[6] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_6__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_5__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_152), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[5] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_5__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_4__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_167), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[4] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_4__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_3__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_182), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[3] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_3__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_2__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_197), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[2] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_2__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_1__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_212), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[1] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_1__i0_i15.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_0__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_227), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[0] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_0__i0_i15.GSR = "ENABLED";
    FD1P3AX address_i0_i1 (.D(cpu_fpga_bus_a_c_1), .SP(cpu_fpga_clk_c_enable_230), 
            .CK(cpu_fpga_clk_c), .Q(address[1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam address_i0_i1.GSR = "ENABLED";
    FD1P3AX address_i0_i2 (.D(cpu_fpga_bus_a_c_2), .SP(cpu_fpga_clk_c_enable_230), 
            .CK(cpu_fpga_clk_c), .Q(address[2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam address_i0_i2.GSR = "ENABLED";
    FD1P3AX address_i0_i3 (.D(cpu_fpga_bus_a_c_3), .SP(cpu_fpga_clk_c_enable_230), 
            .CK(cpu_fpga_clk_c), .Q(address[3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam address_i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i1.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_15__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_245), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[15] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_15__i0_i15.GSR = "ENABLED";
    FD1S3JX STATE_FSM_i2 (.D(n26), .CK(cpu_fpga_clk_c), .PD(n3534), .Q(n1792));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(50[4] 87[13])
    defparam STATE_FSM_i2.GSR = "ENABLED";
    LUT4 i1181_3_lut (.A(\BUFF[8] [6]), .B(\BUFF[9] [6]), .C(\BUFF[0] [0]), 
         .Z(n3121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1181_3_lut.init = 16'hcaca;
    LUT4 i1180_3_lut (.A(\BUFF[6] [6]), .B(\BUFF[7] [6]), .C(\BUFF[0] [0]), 
         .Z(n3120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1180_3_lut.init = 16'hcaca;
    LUT4 i1033_3_lut (.A(\BUFF[12] [8]), .B(\BUFF[13] [8]), .C(address[0]), 
         .Z(n2973)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1033_3_lut.init = 16'hcaca;
    LUT4 i1210_3_lut (.A(\BUFF[6] [1]), .B(\BUFF[7] [1]), .C(\BUFF[0] [0]), 
         .Z(n3150)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1210_3_lut.init = 16'hcaca;
    LUT4 i968_3_lut (.A(\BUFF[2] [2]), .B(\BUFF[3] [2]), .C(\BUFF[0] [0]), 
         .Z(n2908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i968_3_lut.init = 16'hcaca;
    LUT4 i648_1_lut (.A(cpu_fpga_bus_d_15__N_17), .Z(n2626)) /* synthesis lut_function=(!(A)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(33[2] 89[14])
    defparam i648_1_lut.init = 16'h5555;
    LUT4 equal_343_i5_2_lut (.A(address[0]), .B(address[1]), .Z(n5_adj_1)) /* synthesis lut_function=(A+(B)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(70[12:41])
    defparam equal_343_i5_2_lut.init = 16'heeee;
    LUT4 i878_2_lut (.A(address[0]), .B(address[1]), .Z(n2692)) /* synthesis lut_function=(A (B)) */ ;
    defparam i878_2_lut.init = 16'h8888;
    LUT4 i1209_3_lut (.A(\BUFF[4] [1]), .B(\BUFF[5] [1]), .C(\BUFF[0] [0]), 
         .Z(n3149)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1209_3_lut.init = 16'hcaca;
    LUT4 i1139_3_lut (.A(\BUFF[14] [2]), .B(\BUFF[15] [2]), .C(address[0]), 
         .Z(n3079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1139_3_lut.init = 16'hcaca;
    LUT4 i1138_3_lut (.A(\BUFF[12] [2]), .B(\BUFF[13] [2]), .C(address[0]), 
         .Z(n3078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1138_3_lut.init = 16'hcaca;
    LUT4 i1137_3_lut (.A(\BUFF[10] [2]), .B(\BUFF[11] [2]), .C(address[0]), 
         .Z(n3077)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1137_3_lut.init = 16'hcaca;
    LUT4 i1136_3_lut (.A(\BUFF[8] [2]), .B(\BUFF[9] [2]), .C(address[0]), 
         .Z(n3076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1136_3_lut.init = 16'hcaca;
    LUT4 i1135_3_lut (.A(\BUFF[6] [2]), .B(\BUFF[7] [2]), .C(address[0]), 
         .Z(n3075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1135_3_lut.init = 16'hcaca;
    LUT4 i1134_3_lut (.A(\BUFF[4] [2]), .B(\BUFF[5] [2]), .C(address[0]), 
         .Z(n3074)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1134_3_lut.init = 16'hcaca;
    LUT4 i985_3_lut (.A(\BUFF[6] [11]), .B(\BUFF[7] [11]), .C(address[0]), 
         .Z(n2925)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i985_3_lut.init = 16'hcaca;
    LUT4 i984_3_lut (.A(\BUFF[4] [11]), .B(\BUFF[5] [11]), .C(address[0]), 
         .Z(n2924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i984_3_lut.init = 16'hcaca;
    LUT4 i983_3_lut (.A(\BUFF[2] [11]), .B(\BUFF[3] [11]), .C(address[0]), 
         .Z(n2923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i983_3_lut.init = 16'hcaca;
    LUT4 i982_3_lut (.A(\BUFF[0] [11]), .B(\BUFF[1] [11]), .C(address[0]), 
         .Z(n2922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i982_3_lut.init = 16'hcaca;
    LUT4 i1133_3_lut (.A(\BUFF[2] [2]), .B(\BUFF[3] [2]), .C(address[0]), 
         .Z(n3073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1133_3_lut.init = 16'hcaca;
    LUT4 i1132_3_lut (.A(\BUFF[0] [2]), .B(\BUFF[1] [2]), .C(address[0]), 
         .Z(n3072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1132_3_lut.init = 16'hcaca;
    LUT4 i1124_3_lut (.A(\BUFF[14] [3]), .B(\BUFF[15] [3]), .C(address[0]), 
         .Z(n3064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1124_3_lut.init = 16'hcaca;
    LUT4 i1032_3_lut (.A(\BUFF[10] [8]), .B(\BUFF[11] [8]), .C(address[0]), 
         .Z(n2972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1032_3_lut.init = 16'hcaca;
    LUT4 i1123_3_lut (.A(\BUFF[12] [3]), .B(\BUFF[13] [3]), .C(address[0]), 
         .Z(n3063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1123_3_lut.init = 16'hcaca;
    LUT4 i1122_3_lut (.A(\BUFF[10] [3]), .B(\BUFF[11] [3]), .C(address[0]), 
         .Z(n3062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1122_3_lut.init = 16'hcaca;
    LUT4 i1121_3_lut (.A(\BUFF[8] [3]), .B(\BUFF[9] [3]), .C(address[0]), 
         .Z(n3061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1121_3_lut.init = 16'hcaca;
    LUT4 i1120_3_lut (.A(\BUFF[6] [3]), .B(\BUFF[7] [3]), .C(address[0]), 
         .Z(n3060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1120_3_lut.init = 16'hcaca;
    LUT4 i1119_3_lut (.A(\BUFF[4] [3]), .B(\BUFF[5] [3]), .C(address[0]), 
         .Z(n3059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1119_3_lut.init = 16'hcaca;
    LUT4 i1118_3_lut (.A(\BUFF[2] [3]), .B(\BUFF[3] [3]), .C(address[0]), 
         .Z(n3058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1118_3_lut.init = 16'hcaca;
    LUT4 i1117_3_lut (.A(\BUFF[0] [3]), .B(\BUFF[1] [3]), .C(address[0]), 
         .Z(n3057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1117_3_lut.init = 16'hcaca;
    LUT4 i1259_3_lut (.A(\BUFF[14] [13]), .B(\BUFF[15] [13]), .C(address[0]), 
         .Z(n3199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1259_3_lut.init = 16'hcaca;
    LUT4 i1258_3_lut (.A(\BUFF[12] [13]), .B(\BUFF[13] [13]), .C(address[0]), 
         .Z(n3198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1258_3_lut.init = 16'hcaca;
    LUT4 i1257_3_lut (.A(\BUFF[10] [13]), .B(\BUFF[11] [13]), .C(address[0]), 
         .Z(n3197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1257_3_lut.init = 16'hcaca;
    LUT4 i1256_3_lut (.A(\BUFF[8] [13]), .B(\BUFF[9] [13]), .C(address[0]), 
         .Z(n3196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1256_3_lut.init = 16'hcaca;
    LUT4 i1255_3_lut (.A(\BUFF[6] [13]), .B(\BUFF[7] [13]), .C(address[0]), 
         .Z(n3195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1255_3_lut.init = 16'hcaca;
    LUT4 i1254_3_lut (.A(\BUFF[4] [13]), .B(\BUFF[5] [13]), .C(address[0]), 
         .Z(n3194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1254_3_lut.init = 16'hcaca;
    LUT4 i1031_3_lut (.A(\BUFF[8] [8]), .B(\BUFF[9] [8]), .C(address[0]), 
         .Z(n2971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1031_3_lut.init = 16'hcaca;
    LUT4 i1319_3_lut (.A(\BUFF[14] [3]), .B(\BUFF[15] [3]), .C(\BUFF[0] [0]), 
         .Z(n3259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1319_3_lut.init = 16'hcaca;
    LUT4 i1318_3_lut (.A(\BUFF[12] [3]), .B(\BUFF[13] [3]), .C(\BUFF[0] [0]), 
         .Z(n3258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1318_3_lut.init = 16'hcaca;
    LUT4 i1253_3_lut (.A(\BUFF[2] [13]), .B(\BUFF[3] [13]), .C(address[0]), 
         .Z(n3193)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1253_3_lut.init = 16'hcaca;
    LUT4 i1252_3_lut (.A(\BUFF[0] [13]), .B(\BUFF[1] [13]), .C(address[0]), 
         .Z(n3192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1252_3_lut.init = 16'hcaca;
    LUT4 i1109_3_lut (.A(\BUFF[14] [4]), .B(\BUFF[15] [4]), .C(address[0]), 
         .Z(n3049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1109_3_lut.init = 16'hcaca;
    LUT4 i1108_3_lut (.A(\BUFF[12] [4]), .B(\BUFF[13] [4]), .C(address[0]), 
         .Z(n3048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1108_3_lut.init = 16'hcaca;
    LUT4 i1317_3_lut (.A(\BUFF[10] [3]), .B(\BUFF[11] [3]), .C(\BUFF[0] [0]), 
         .Z(n3257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1317_3_lut.init = 16'hcaca;
    LUT4 i1316_3_lut (.A(\BUFF[8] [3]), .B(\BUFF[9] [3]), .C(\BUFF[0] [0]), 
         .Z(n3256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1316_3_lut.init = 16'hcaca;
    LUT4 i1107_3_lut (.A(\BUFF[10] [4]), .B(\BUFF[11] [4]), .C(address[0]), 
         .Z(n3047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1107_3_lut.init = 16'hcaca;
    LUT4 i1106_3_lut (.A(\BUFF[8] [4]), .B(\BUFF[9] [4]), .C(address[0]), 
         .Z(n3046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1106_3_lut.init = 16'hcaca;
    LUT4 i1105_3_lut (.A(\BUFF[6] [4]), .B(\BUFF[7] [4]), .C(address[0]), 
         .Z(n3045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1105_3_lut.init = 16'hcaca;
    LUT4 i1104_3_lut (.A(\BUFF[4] [4]), .B(\BUFF[5] [4]), .C(address[0]), 
         .Z(n3044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1104_3_lut.init = 16'hcaca;
    LUT4 i1103_3_lut (.A(\BUFF[2] [4]), .B(\BUFF[3] [4]), .C(address[0]), 
         .Z(n3043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1103_3_lut.init = 16'hcaca;
    LUT4 i1030_3_lut (.A(\BUFF[6] [8]), .B(\BUFF[7] [8]), .C(address[0]), 
         .Z(n2970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1030_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n3534), .B(address[3]), .C(n2692), .D(address[2]), 
         .Z(cpu_fpga_clk_c_enable_182)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1 (.A(n3534), .B(address[3]), .C(n5_adj_2), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_197)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_4_lut_adj_2 (.A(n3534), .B(address[3]), .C(n5), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_212)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_2.init = 16'h0002;
    LUT4 i1102_3_lut (.A(\BUFF[0] [4]), .B(\BUFF[1] [4]), .C(address[0]), 
         .Z(n3042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1102_3_lut.init = 16'hcaca;
    LUT4 i1315_3_lut (.A(\BUFF[6] [3]), .B(\BUFF[7] [3]), .C(\BUFF[0] [0]), 
         .Z(n3255)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1315_3_lut.init = 16'hcaca;
    LUT4 i1314_3_lut (.A(\BUFF[4] [3]), .B(\BUFF[5] [3]), .C(\BUFF[0] [0]), 
         .Z(n3254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1314_3_lut.init = 16'hcaca;
    LUT4 i1313_3_lut (.A(\BUFF[2] [3]), .B(\BUFF[3] [3]), .C(\BUFF[0] [0]), 
         .Z(n3253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1313_3_lut.init = 16'hcaca;
    LUT4 i1091_3_lut (.A(\BUFF[8] [0]), .B(\BUFF[9] [0]), .C(address[0]), 
         .Z(n3031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1091_3_lut.init = 16'hcaca;
    LUT4 i1090_3_lut (.A(\BUFF[6] [0]), .B(\BUFF[7] [0]), .C(address[0]), 
         .Z(n3030)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1090_3_lut.init = 16'hcaca;
    LUT4 i1089_3_lut (.A(\BUFF[4] [0]), .B(\BUFF[5] [0]), .C(address[0]), 
         .Z(n3029)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1089_3_lut.init = 16'hcaca;
    LUT4 i1088_3_lut (.A(\BUFF[2] [0]), .B(\BUFF[3] [0]), .C(address[0]), 
         .Z(n3028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1088_3_lut.init = 16'hcaca;
    LUT4 i1087_3_lut (.A(\BUFF[0] [0]), .B(\BUFF[1] [0]), .C(address[0]), 
         .Z(n3027)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1087_3_lut.init = 16'hcaca;
    LUT4 i1244_3_lut (.A(\BUFF[14] [14]), .B(\BUFF[15] [14]), .C(address[0]), 
         .Z(n3184)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1244_3_lut.init = 16'hcaca;
    LUT4 i1029_3_lut (.A(\BUFF[4] [8]), .B(\BUFF[5] [8]), .C(address[0]), 
         .Z(n2969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1029_3_lut.init = 16'hcaca;
    LUT4 i1243_3_lut (.A(\BUFF[12] [14]), .B(\BUFF[13] [14]), .C(address[0]), 
         .Z(n3183)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1243_3_lut.init = 16'hcaca;
    LUT4 i1242_3_lut (.A(\BUFF[10] [14]), .B(\BUFF[11] [14]), .C(address[0]), 
         .Z(n3182)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1242_3_lut.init = 16'hcaca;
    LUT4 i1241_3_lut (.A(\BUFF[8] [14]), .B(\BUFF[9] [14]), .C(address[0]), 
         .Z(n3181)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1241_3_lut.init = 16'hcaca;
    LUT4 i1240_3_lut (.A(\BUFF[6] [14]), .B(\BUFF[7] [14]), .C(address[0]), 
         .Z(n3180)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1240_3_lut.init = 16'hcaca;
    LUT4 i1239_3_lut (.A(\BUFF[4] [14]), .B(\BUFF[5] [14]), .C(address[0]), 
         .Z(n3179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1239_3_lut.init = 16'hcaca;
    LUT4 i1238_3_lut (.A(\BUFF[2] [14]), .B(\BUFF[3] [14]), .C(address[0]), 
         .Z(n3178)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1238_3_lut.init = 16'hcaca;
    LUT4 i1237_3_lut (.A(\BUFF[0] [14]), .B(\BUFF[1] [14]), .C(address[0]), 
         .Z(n3177)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1237_3_lut.init = 16'hcaca;
    LUT4 i1079_3_lut (.A(\BUFF[14] [5]), .B(\BUFF[15] [5]), .C(address[0]), 
         .Z(n3019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1079_3_lut.init = 16'hcaca;
    LUT4 i1078_3_lut (.A(\BUFF[12] [5]), .B(\BUFF[13] [5]), .C(address[0]), 
         .Z(n3018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1078_3_lut.init = 16'hcaca;
    L6MUX21 i1971 (.D0(n3777), .D1(n3774), .SD(address[2]), .Z(n3778));
    LUT4 i1208_3_lut (.A(\BUFF[2] [1]), .B(\BUFF[3] [1]), .C(\BUFF[0] [0]), 
         .Z(n3148)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1208_3_lut.init = 16'hcaca;
    PFUMX i1969 (.BLUT(n3776), .ALUT(n3775), .C0(address[0]), .Z(n3777));
    LUT4 i1207_3_lut (.A(\BUFF[0] [1]), .B(\BUFF[1] [1]), .C(\BUFF[0] [0]), 
         .Z(n3147)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1207_3_lut.init = 16'hcaca;
    LUT4 i967_3_lut (.A(\BUFF[0] [2]), .B(\BUFF[1] [2]), .C(\BUFF[0] [0]), 
         .Z(n2907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i967_3_lut.init = 16'hcaca;
    PFUMX i1966 (.BLUT(n3773), .ALUT(n3772), .C0(address[0]), .Z(n3774));
    LUT4 i1028_3_lut (.A(\BUFF[2] [8]), .B(\BUFF[3] [8]), .C(address[0]), 
         .Z(n2968)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1028_3_lut.init = 16'hcaca;
    L6MUX21 i1963 (.D0(n3770), .D1(n3767), .SD(address[2]), .Z(n3771));
    LUT4 i1027_3_lut (.A(\BUFF[0] [8]), .B(\BUFF[1] [8]), .C(address[0]), 
         .Z(n2967)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1027_3_lut.init = 16'hcaca;
    PFUMX i1961 (.BLUT(n3769), .ALUT(n3768), .C0(address[0]), .Z(n3770));
    LUT4 i1019_3_lut (.A(\BUFF[14] [9]), .B(\BUFF[15] [9]), .C(address[0]), 
         .Z(n2959)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1019_3_lut.init = 16'hcaca;
    PFUMX i1958 (.BLUT(n3766), .ALUT(n3765), .C0(address[0]), .Z(n3767));
    LUT4 i1179_3_lut (.A(\BUFF[4] [6]), .B(\BUFF[5] [6]), .C(\BUFF[0] [0]), 
         .Z(n3119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1179_3_lut.init = 16'hcaca;
    LUT4 i1018_3_lut (.A(\BUFF[12] [9]), .B(\BUFF[13] [9]), .C(address[0]), 
         .Z(n2958)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1018_3_lut.init = 16'hcaca;
    L6MUX21 i1955 (.D0(n3763), .D1(n3760), .SD(address[2]), .Z(n3764));
    LUT4 i1017_3_lut (.A(\BUFF[10] [9]), .B(\BUFF[11] [9]), .C(address[0]), 
         .Z(n2957)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1017_3_lut.init = 16'hcaca;
    PFUMX i1953 (.BLUT(n3762), .ALUT(n3761), .C0(address[0]), .Z(n3763));
    LUT4 i1016_3_lut (.A(\BUFF[8] [9]), .B(\BUFF[9] [9]), .C(address[0]), 
         .Z(n2956)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1016_3_lut.init = 16'hcaca;
    PFUMX i1950 (.BLUT(n3759), .ALUT(n3758), .C0(address[0]), .Z(n3760));
    LUT4 i1015_3_lut (.A(\BUFF[6] [9]), .B(\BUFF[7] [9]), .C(address[0]), 
         .Z(n2955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1015_3_lut.init = 16'hcaca;
    PFUMX i1170 (.BLUT(n3102), .ALUT(n3103), .C0(\BUFF[0] [1]), .Z(n3110));
    L6MUX21 i1947 (.D0(n3756), .D1(n3753), .SD(address[2]), .Z(n3757));
    LUT4 i1014_3_lut (.A(\BUFF[4] [9]), .B(\BUFF[5] [9]), .C(address[0]), 
         .Z(n2954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1014_3_lut.init = 16'hcaca;
    PFUMX i1945 (.BLUT(n3755), .ALUT(n3754), .C0(address[0]), .Z(n3756));
    LUT4 i1013_3_lut (.A(\BUFF[2] [9]), .B(\BUFF[3] [9]), .C(address[0]), 
         .Z(n2953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1013_3_lut.init = 16'hcaca;
    PFUMX i1942 (.BLUT(n3752), .ALUT(n3751), .C0(address[0]), .Z(n3753));
    LUT4 i1012_3_lut (.A(\BUFF[0] [9]), .B(\BUFF[1] [9]), .C(address[0]), 
         .Z(n2952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1012_3_lut.init = 16'hcaca;
    LUT4 i1199_3_lut (.A(\BUFF[14] [5]), .B(\BUFF[15] [5]), .C(\BUFF[0] [0]), 
         .Z(n3139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1199_3_lut.init = 16'hcaca;
    LUT4 i1198_3_lut (.A(\BUFF[12] [5]), .B(\BUFF[13] [5]), .C(\BUFF[0] [0]), 
         .Z(n3138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1198_3_lut.init = 16'hcaca;
    LUT4 i1197_3_lut (.A(\BUFF[10] [5]), .B(\BUFF[11] [5]), .C(\BUFF[0] [0]), 
         .Z(n3137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1197_3_lut.init = 16'hcaca;
    LUT4 i1196_3_lut (.A(\BUFF[8] [5]), .B(\BUFF[9] [5]), .C(\BUFF[0] [0]), 
         .Z(n3136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1196_3_lut.init = 16'hcaca;
    LUT4 i1195_3_lut (.A(\BUFF[6] [5]), .B(\BUFF[7] [5]), .C(\BUFF[0] [0]), 
         .Z(n3135)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1195_3_lut.init = 16'hcaca;
    LUT4 i1194_3_lut (.A(\BUFF[4] [5]), .B(\BUFF[5] [5]), .C(\BUFF[0] [0]), 
         .Z(n3134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1194_3_lut.init = 16'hcaca;
    LUT4 i1289_3_lut (.A(\BUFF[14] [7]), .B(\BUFF[15] [7]), .C(\BUFF[0] [0]), 
         .Z(n3229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1289_3_lut.init = 16'hcaca;
    LUT4 i1288_3_lut (.A(\BUFF[12] [7]), .B(\BUFF[13] [7]), .C(\BUFF[0] [0]), 
         .Z(n3228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1288_3_lut.init = 16'hcaca;
    LUT4 i1193_3_lut (.A(\BUFF[2] [5]), .B(\BUFF[3] [5]), .C(\BUFF[0] [0]), 
         .Z(n3133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1193_3_lut.init = 16'hcaca;
    LUT4 i1192_3_lut (.A(\BUFF[0] [5]), .B(\BUFF[1] [5]), .C(\BUFF[0] [0]), 
         .Z(n3132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1192_3_lut.init = 16'hcaca;
    LUT4 i1004_3_lut (.A(\BUFF[14] [10]), .B(\BUFF[15] [10]), .C(address[0]), 
         .Z(n2944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1004_3_lut.init = 16'hcaca;
    LUT4 i1003_3_lut (.A(\BUFF[12] [10]), .B(\BUFF[13] [10]), .C(address[0]), 
         .Z(n2943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1003_3_lut.init = 16'hcaca;
    LUT4 i1287_3_lut (.A(\BUFF[10] [7]), .B(\BUFF[11] [7]), .C(\BUFF[0] [0]), 
         .Z(n3227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1287_3_lut.init = 16'hcaca;
    LUT4 i1286_3_lut (.A(\BUFF[8] [7]), .B(\BUFF[9] [7]), .C(\BUFF[0] [0]), 
         .Z(n3226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1286_3_lut.init = 16'hcaca;
    LUT4 i1002_3_lut (.A(\BUFF[10] [10]), .B(\BUFF[11] [10]), .C(address[0]), 
         .Z(n2942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1002_3_lut.init = 16'hcaca;
    LUT4 i1001_3_lut (.A(\BUFF[8] [10]), .B(\BUFF[9] [10]), .C(address[0]), 
         .Z(n2941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1001_3_lut.init = 16'hcaca;
    LUT4 i1000_3_lut (.A(\BUFF[6] [10]), .B(\BUFF[7] [10]), .C(address[0]), 
         .Z(n2940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1000_3_lut.init = 16'hcaca;
    LUT4 i999_3_lut (.A(\BUFF[4] [10]), .B(\BUFF[5] [10]), .C(address[0]), 
         .Z(n2939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i999_3_lut.init = 16'hcaca;
    LUT4 i998_3_lut (.A(\BUFF[2] [10]), .B(\BUFF[3] [10]), .C(address[0]), 
         .Z(n2938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i998_3_lut.init = 16'hcaca;
    LUT4 i997_3_lut (.A(\BUFF[0] [10]), .B(\BUFF[1] [10]), .C(address[0]), 
         .Z(n2937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i997_3_lut.init = 16'hcaca;
    LUT4 i1285_3_lut (.A(\BUFF[6] [7]), .B(\BUFF[7] [7]), .C(\BUFF[0] [0]), 
         .Z(n3225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1285_3_lut.init = 16'hcaca;
    LUT4 i1284_3_lut (.A(\BUFF[4] [7]), .B(\BUFF[5] [7]), .C(\BUFF[0] [0]), 
         .Z(n3224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1284_3_lut.init = 16'hcaca;
    LUT4 i1283_3_lut (.A(\BUFF[2] [7]), .B(\BUFF[3] [7]), .C(\BUFF[0] [0]), 
         .Z(n3223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1283_3_lut.init = 16'hcaca;
    LUT4 i1282_3_lut (.A(\BUFF[0] [7]), .B(\BUFF[1] [7]), .C(\BUFF[0] [0]), 
         .Z(n3222)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1282_3_lut.init = 16'hcaca;
    LUT4 i1184_3_lut (.A(\BUFF[14] [6]), .B(\BUFF[15] [6]), .C(\BUFF[0] [0]), 
         .Z(n3124)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1184_3_lut.init = 16'hcaca;
    LUT4 i1165_3_lut (.A(\BUFF[6] [0]), .B(\BUFF[7] [0]), .C(\BUFF[0] [0]), 
         .Z(n3105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1165_3_lut.init = 16'hcaca;
    LUT4 equal_337_i5_2_lut (.A(address[0]), .B(address[1]), .Z(n5_adj_2)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(70[12:41])
    defparam equal_337_i5_2_lut.init = 16'hbbbb;
    LUT4 equal_342_i5_2_lut (.A(address[0]), .B(address[1]), .Z(n5)) /* synthesis lut_function=((B)+!A) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(70[12:41])
    defparam equal_342_i5_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut_adj_3 (.A(n3534), .B(address[3]), .C(n5_adj_1), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_227)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_3.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_4_lut_adj_4 (.A(n3534), .B(address[3]), .C(n2692), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_122)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_4.init = 16'h2000;
    FD1S3AX STATE_FSM_i3 (.D(n2655), .CK(cpu_fpga_clk_c), .Q(n1791));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(50[4] 87[13])
    defparam STATE_FSM_i3.GSR = "ENABLED";
    FD1S3AX STATE_FSM_i4 (.D(n2661), .CK(cpu_fpga_clk_c), .Q(n1790));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(50[4] 87[13])
    defparam STATE_FSM_i4.GSR = "ENABLED";
    FD1S3AX STATE_FSM_i5 (.D(n13), .CK(cpu_fpga_clk_c), .Q(n1789));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(50[4] 87[13])
    defparam STATE_FSM_i5.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i1 (.D(cpu_fpga_bus_d_15__N_570[1]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i1.GSR = "ENABLED";
    LUT4 i1164_3_lut (.A(\BUFF[4] [0]), .B(\BUFF[5] [0]), .C(\BUFF[0] [0]), 
         .Z(n3104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1164_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_5 (.A(n3534), .B(address[3]), .C(n5_adj_2), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_137)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_5.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_6 (.A(n3534), .B(address[3]), .C(n5), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_152)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_6.init = 16'h0200;
    LUT4 i1_3_lut (.A(STATE_2__N_297_c_0), .B(n1791), .C(cpu_fpga_bus_nwe_c), 
         .Z(cpu_fpga_clk_c_enable_230)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B))) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(23[9:14])
    defparam i1_3_lut.init = 16'h4c4c;
    LUT4 i769_1_lut (.A(cpu_fpga_rst_c), .Z(n2760)) /* synthesis lut_function=(!(A)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(14[4:16])
    defparam i769_1_lut.init = 16'h5555;
    LUT4 fpga_io_gp_7__I_0_i1_1_lut (.A(fpga_io_gp_7__N_18[0]), .Z(fpga_io_gp_c_0)) /* synthesis lut_function=(!(A)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(91[20:55])
    defparam fpga_io_gp_7__I_0_i1_1_lut.init = 16'h5555;
    LUT4 fpga_io_gp_7__I_0_i2_1_lut (.A(fpga_io_gp_7__N_18[1]), .Z(fpga_io_gp_c_1)) /* synthesis lut_function=(!(A)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(91[20:55])
    defparam fpga_io_gp_7__I_0_i2_1_lut.init = 16'h5555;
    LUT4 fpga_io_gp_7__I_0_i3_1_lut (.A(fpga_io_gp_7__N_18[2]), .Z(fpga_io_gp_c_2)) /* synthesis lut_function=(!(A)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(91[20:55])
    defparam fpga_io_gp_7__I_0_i3_1_lut.init = 16'h5555;
    LUT4 fpga_io_gp_7__I_0_i4_1_lut (.A(fpga_io_gp_7__N_18[3]), .Z(fpga_io_gp_c_3)) /* synthesis lut_function=(!(A)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(91[20:55])
    defparam fpga_io_gp_7__I_0_i4_1_lut.init = 16'h5555;
    LUT4 fpga_io_gp_7__I_0_i5_1_lut (.A(fpga_io_gp_7__N_18[4]), .Z(fpga_io_gp_c_4)) /* synthesis lut_function=(!(A)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(91[20:55])
    defparam fpga_io_gp_7__I_0_i5_1_lut.init = 16'h5555;
    LUT4 i770_1_lut (.A(n1789), .Z(n2761)) /* synthesis lut_function=(!(A)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(50[4] 87[13])
    defparam i770_1_lut.init = 16'h5555;
    LUT4 fpga_io_gp_7__I_0_i6_1_lut (.A(fpga_io_gp_7__N_18[5]), .Z(fpga_io_gp_c_5)) /* synthesis lut_function=(!(A)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(91[20:55])
    defparam fpga_io_gp_7__I_0_i6_1_lut.init = 16'h5555;
    LUT4 fpga_io_gp_7__I_0_i7_1_lut (.A(fpga_io_gp_7__N_18[6]), .Z(fpga_io_gp_c_6)) /* synthesis lut_function=(!(A)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(91[20:55])
    defparam fpga_io_gp_7__I_0_i7_1_lut.init = 16'h5555;
    LUT4 fpga_io_gp_7__I_0_i8_1_lut (.A(fpga_io_gp_7__N_18[7]), .Z(fpga_io_gp_c_7)) /* synthesis lut_function=(!(A)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(91[20:55])
    defparam fpga_io_gp_7__I_0_i8_1_lut.init = 16'h5555;
    LUT4 i1_4_lut (.A(STATE_2__N_297_c_0), .B(n1792), .C(n1789), .D(cpu_fpga_bus_ne1_c), 
         .Z(n26)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(23[9:14])
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i1_4_lut_adj_7 (.A(STATE_2__N_297_c_0), .B(n1792), .C(n3532), 
         .D(cpu_fpga_bus_ne1_c), .Z(n2655)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(23[9:14])
    defparam i1_4_lut_adj_7.init = 16'ha0ec;
    PFUMX i1171 (.BLUT(n3104), .ALUT(n3105), .C0(\BUFF[0] [1]), .Z(n3111));
    LUT4 i1_3_lut_adj_8 (.A(cpu_fpga_bus_nwe_c), .B(n1790), .C(n1791), 
         .Z(n2661)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(10[4:20])
    defparam i1_3_lut_adj_8.init = 16'h5454;
    LUT4 i1_2_lut_3_lut_4_lut_adj_9 (.A(n3534), .B(address[3]), .C(n5_adj_1), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_167)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_9.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_10 (.A(address[3]), .B(n3534), .C(n5_adj_2), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_77)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_10.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_11 (.A(address[3]), .B(n3534), .C(n2692), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_62)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_11.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_12 (.A(address[3]), .B(n3534), .C(n5), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_92)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_12.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_13 (.A(address[3]), .B(n3534), .C(n5_adj_1), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_107)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_13.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_14 (.A(address[3]), .B(n3534), .C(n5_adj_1), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_47)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_14.init = 16'h0800;
    LUT4 i1094_3_lut (.A(\BUFF[14] [0]), .B(\BUFF[15] [0]), .C(address[0]), 
         .Z(n3034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1094_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_15 (.A(address[3]), .B(n3534), .C(n2692), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_245)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_15.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_16 (.A(address[3]), .B(n3534), .C(n5), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_32)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_16.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_17 (.A(address[3]), .B(n3534), .C(n5_adj_2), 
         .D(address[2]), .Z(cpu_fpga_clk_c_enable_260)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_17.init = 16'h0800;
    LUT4 i1_2_lut_rep_11 (.A(n1791), .B(cpu_fpga_bus_nwe_c), .Z(n3532)) /* synthesis lut_function=(A (B)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(50[4] 87[13])
    defparam i1_2_lut_rep_11.init = 16'h8888;
    LUT4 cpu_fpga_bus_noe_I_0_1_lut_rep_12 (.A(STATE_2__N_297_c_0), .Z(n3533)) /* synthesis lut_function=(!(A)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(61[12:34])
    defparam cpu_fpga_bus_noe_I_0_1_lut_rep_12.init = 16'h5555;
    LUT4 i1_3_lut_4_lut_4_lut (.A(STATE_2__N_297_c_0), .B(n1789), .C(cpu_fpga_bus_nwe_c), 
         .D(n1791), .Z(n13)) /* synthesis lut_function=(!(A+!(B+(C (D))))) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(61[12:34])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h5444;
    LUT4 i1_2_lut_rep_13 (.A(cpu_fpga_bus_nwe_c), .B(n1790), .Z(n3534)) /* synthesis lut_function=(A (B)) */ ;   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(10[4:20])
    defparam i1_2_lut_rep_13.init = 16'h8888;
    LUT4 i1163_3_lut (.A(\BUFF[2] [0]), .B(\BUFF[3] [0]), .C(\BUFF[0] [0]), 
         .Z(n3103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1163_3_lut.init = 16'hcaca;
    MUX21 i1526 (.D0(n2949), .D1(n2950), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[10]));
    LUT4 \BUFF_13[[12__bdd_3_lut  (.A(\BUFF[12] [12]), .B(\BUFF[14] [12]), 
         .C(address[1]), .Z(n3752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_13[[12__bdd_3_lut .init = 16'hcaca;
    PFUMX i1290 (.BLUT(n3222), .ALUT(n3223), .C0(\BUFF[0] [1]), .Z(n3230));
    PFUMX i1291 (.BLUT(n3224), .ALUT(n3225), .C0(\BUFF[0] [1]), .Z(n3231));
    PFUMX i1005 (.BLUT(n2937), .ALUT(n2938), .C0(address[1]), .Z(n2945));
    PFUMX i1006 (.BLUT(n2939), .ALUT(n2940), .C0(address[1]), .Z(n2946));
    PFUMX i1007 (.BLUT(n2941), .ALUT(n2942), .C0(address[1]), .Z(n2947));
    PFUMX i1292 (.BLUT(n3226), .ALUT(n3227), .C0(\BUFF[0] [1]), .Z(n3232));
    PFUMX i1008 (.BLUT(n2943), .ALUT(n2944), .C0(address[1]), .Z(n2948));
    PFUMX i1200 (.BLUT(n3132), .ALUT(n3133), .C0(\BUFF[0] [1]), .Z(n3140));
    PFUMX i1293 (.BLUT(n3228), .ALUT(n3229), .C0(\BUFF[0] [1]), .Z(n3233));
    PFUMX i1201 (.BLUT(n3134), .ALUT(n3135), .C0(\BUFF[0] [1]), .Z(n3141));
    PFUMX i1202 (.BLUT(n3136), .ALUT(n3137), .C0(\BUFF[0] [1]), .Z(n3142));
    PFUMX i1203 (.BLUT(n3138), .ALUT(n3139), .C0(\BUFF[0] [1]), .Z(n3143));
    PFUMX i1020 (.BLUT(n2952), .ALUT(n2953), .C0(address[1]), .Z(n2960));
    PFUMX i1021 (.BLUT(n2954), .ALUT(n2955), .C0(address[1]), .Z(n2961));
    PFUMX i1022 (.BLUT(n2956), .ALUT(n2957), .C0(address[1]), .Z(n2962));
    PFUMX i1023 (.BLUT(n2958), .ALUT(n2959), .C0(address[1]), .Z(n2963));
    PFUMX i1035 (.BLUT(n2967), .ALUT(n2968), .C0(address[1]), .Z(n2975));
    PFUMX i1215 (.BLUT(n3147), .ALUT(n3148), .C0(\BUFF[0] [1]), .Z(n3155));
    PFUMX i1036 (.BLUT(n2969), .ALUT(n2970), .C0(address[1]), .Z(n2976));
    PFUMX i1037 (.BLUT(n2971), .ALUT(n2972), .C0(address[1]), .Z(n2977));
    PFUMX i1216 (.BLUT(n3149), .ALUT(n3150), .C0(\BUFF[0] [1]), .Z(n3156));
    PFUMX i1038 (.BLUT(n2973), .ALUT(n2974), .C0(address[1]), .Z(n2978));
    PFUMX i1217 (.BLUT(n3151), .ALUT(n3152), .C0(\BUFF[0] [1]), .Z(n3157));
    PFUMX i1218 (.BLUT(n3153), .ALUT(n3154), .C0(\BUFF[0] [1]), .Z(n3158));
    PFUMX i1050 (.BLUT(n2982), .ALUT(n2983), .C0(address[1]), .Z(n2990));
    PFUMX i1051 (.BLUT(n2984), .ALUT(n2985), .C0(address[1]), .Z(n2991));
    PFUMX i1052 (.BLUT(n2986), .ALUT(n2987), .C0(address[1]), .Z(n2992));
    PFUMX i1305 (.BLUT(n3237), .ALUT(n3238), .C0(\BUFF[0] [1]), .Z(n3245));
    PFUMX i1053 (.BLUT(n2988), .ALUT(n2989), .C0(address[1]), .Z(n2993));
    PFUMX i1306 (.BLUT(n3239), .ALUT(n3240), .C0(\BUFF[0] [1]), .Z(n3246));
    PFUMX i1307 (.BLUT(n3241), .ALUT(n3242), .C0(\BUFF[0] [1]), .Z(n3247));
    PFUMX i1230 (.BLUT(n3162), .ALUT(n3163), .C0(address[1]), .Z(n3170));
    PFUMX i1308 (.BLUT(n3243), .ALUT(n3244), .C0(\BUFF[0] [1]), .Z(n3248));
    PFUMX i1231 (.BLUT(n3164), .ALUT(n3165), .C0(address[1]), .Z(n3171));
    PFUMX i1065 (.BLUT(n2997), .ALUT(n2998), .C0(address[1]), .Z(n3005));
    PFUMX i1232 (.BLUT(n3166), .ALUT(n3167), .C0(address[1]), .Z(n3172));
    PFUMX i1066 (.BLUT(n2999), .ALUT(n3000), .C0(address[1]), .Z(n3006));
    PFUMX i1067 (.BLUT(n3001), .ALUT(n3002), .C0(address[1]), .Z(n3007));
    PFUMX i1233 (.BLUT(n3168), .ALUT(n3169), .C0(address[1]), .Z(n3173));
    PFUMX i1068 (.BLUT(n3003), .ALUT(n3004), .C0(address[1]), .Z(n3008));
    PFUMX i1080 (.BLUT(n3012), .ALUT(n3013), .C0(address[1]), .Z(n3020));
    FD1S3IX cpu_fpga_bus_d__i2 (.D(cpu_fpga_bus_d_15__N_570[2]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i2.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i3 (.D(cpu_fpga_bus_d_15__N_570[3]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i3.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i4 (.D(cpu_fpga_bus_d_15__N_570[4]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i4.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i5 (.D(cpu_fpga_bus_d_15__N_570[5]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i5.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i6 (.D(cpu_fpga_bus_d_15__N_570[6]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i6.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i7 (.D(cpu_fpga_bus_d_15__N_570[7]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i7.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i8 (.D(cpu_fpga_bus_d_15__N_570[8]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i8.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i9 (.D(cpu_fpga_bus_d_15__N_570[9]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i9.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i10 (.D(cpu_fpga_bus_d_15__N_570[10]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i10.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i11 (.D(cpu_fpga_bus_d_15__N_570[11]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i11.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i12 (.D(cpu_fpga_bus_d_15__N_570[12]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i12.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i13 (.D(cpu_fpga_bus_d_15__N_570[13]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i13.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i14 (.D(cpu_fpga_bus_d_15__N_570[14]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i14.GSR = "ENABLED";
    FD1S3IX cpu_fpga_bus_d__i15 (.D(cpu_fpga_bus_d_15__N_570[15]), .CK(cpu_fpga_clk_c), 
            .CD(n2761), .Q(cpu_fpga_bus_d_15__N_1[15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam cpu_fpga_bus_d__i15.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i1 (.D(cpu_fpga_bus_d_out_1), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [1]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i1.GSR = "ENABLED";
    PFUMX i1081 (.BLUT(n3014), .ALUT(n3015), .C0(address[1]), .Z(n3021));
    PFUMX i1082 (.BLUT(n3016), .ALUT(n3017), .C0(address[1]), .Z(n3022));
    PFUMX i1083 (.BLUT(n3018), .ALUT(n3019), .C0(address[1]), .Z(n3023));
    PFUMX i1245 (.BLUT(n3177), .ALUT(n3178), .C0(address[1]), .Z(n3185));
    PFUMX i1246 (.BLUT(n3179), .ALUT(n3180), .C0(address[1]), .Z(n3186));
    PFUMX i1247 (.BLUT(n3181), .ALUT(n3182), .C0(address[1]), .Z(n3187));
    PFUMX i1248 (.BLUT(n3183), .ALUT(n3184), .C0(address[1]), .Z(n3188));
    PFUMX i1095 (.BLUT(n3027), .ALUT(n3028), .C0(address[1]), .Z(n3035));
    PFUMX i1096 (.BLUT(n3029), .ALUT(n3030), .C0(address[1]), .Z(n3036));
    PFUMX i1321 (.BLUT(n3254), .ALUT(n3255), .C0(\BUFF[0] [1]), .Z(n3261));
    PFUMX i1110 (.BLUT(n3042), .ALUT(n3043), .C0(address[1]), .Z(n3050));
    LUT4 i1162_3_lut (.A(\BUFF[1] [0]), .B(\BUFF[0] [0]), .Z(n3102)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1162_3_lut.init = 16'h8888;
    LUT4 \BUFF_13[[12__bdd_3_lut_1941  (.A(\BUFF[13] [12]), .B(\BUFF[15] [12]), 
         .C(address[1]), .Z(n3751)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_13[[12__bdd_3_lut_1941 .init = 16'hcaca;
    LUT4 \BUFF_8[[12__bdd_3_lut_1944  (.A(\BUFF[11] [12]), .B(\BUFF[9] [12]), 
         .C(address[1]), .Z(n3754)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam \BUFF_8[[12__bdd_3_lut_1944 .init = 16'hacac;
    LUT4 \BUFF_8[[12__bdd_3_lut  (.A(\BUFF[8] [12]), .B(\BUFF[10] [12]), 
         .C(address[1]), .Z(n3755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_8[[12__bdd_3_lut .init = 16'hcaca;
    LUT4 \BUFF_13[[1__bdd_3_lut_1949  (.A(\BUFF[13] [1]), .B(\BUFF[15] [1]), 
         .C(address[1]), .Z(n3758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_13[[1__bdd_3_lut_1949 .init = 16'hcaca;
    LUT4 \BUFF_13[[1__bdd_3_lut  (.A(\BUFF[12] [1]), .B(\BUFF[14] [1]), 
         .C(address[1]), .Z(n3759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_13[[1__bdd_3_lut .init = 16'hcaca;
    LUT4 \BUFF_8[[1__bdd_3_lut_1952  (.A(\BUFF[11] [1]), .B(\BUFF[9] [1]), 
         .C(address[1]), .Z(n3761)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam \BUFF_8[[1__bdd_3_lut_1952 .init = 16'hacac;
    LUT4 i1178_3_lut (.A(\BUFF[2] [6]), .B(\BUFF[3] [6]), .C(\BUFF[0] [0]), 
         .Z(n3118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1178_3_lut.init = 16'hcaca;
    LUT4 \BUFF_8[[1__bdd_3_lut  (.A(\BUFF[8] [1]), .B(\BUFF[10] [1]), .C(address[1]), 
         .Z(n3762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_8[[1__bdd_3_lut .init = 16'hcaca;
    LUT4 i1093_3_lut (.A(\BUFF[12] [0]), .B(\BUFF[13] [0]), .C(address[0]), 
         .Z(n3033)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1093_3_lut.init = 16'hcaca;
    LUT4 i1167_3_lut (.A(\BUFF[10] [0]), .B(\BUFF[11] [0]), .C(\BUFF[0] [0]), 
         .Z(n3107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1167_3_lut.init = 16'hcaca;
    PFUMX i1111 (.BLUT(n3044), .ALUT(n3045), .C0(address[1]), .Z(n3051));
    PFUMX i1112 (.BLUT(n3046), .ALUT(n3047), .C0(address[1]), .Z(n3052));
    MUX21 i1516 (.D0(n3204), .D1(n3205), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[13]));
    LUT4 i1166_3_lut (.A(\BUFF[8] [0]), .B(\BUFF[9] [0]), .C(\BUFF[0] [0]), 
         .Z(n3106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1166_3_lut.init = 16'hcaca;
    LUT4 \BUFF_0[[1__bdd_3_lut_1936  (.A(\BUFF[3] [1]), .B(\BUFF[1] [1]), 
         .C(address[1]), .Z(n3747)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam \BUFF_0[[1__bdd_3_lut_1936 .init = 16'hacac;
    PFUMX i1097 (.BLUT(n3031), .ALUT(n3032), .C0(address[1]), .Z(n3037));
    PFUMX i1322 (.BLUT(n3256), .ALUT(n3257), .C0(\BUFF[0] [1]), .Z(n3262));
    PFUMX i1113 (.BLUT(n3048), .ALUT(n3049), .C0(address[1]), .Z(n3053));
    PFUMX i1260 (.BLUT(n3192), .ALUT(n3193), .C0(address[1]), .Z(n3200));
    PFUMX i1323 (.BLUT(n3258), .ALUT(n3259), .C0(\BUFF[0] [1]), .Z(n3263));
    PFUMX i1261 (.BLUT(n3194), .ALUT(n3195), .C0(address[1]), .Z(n3201));
    PFUMX i1262 (.BLUT(n3196), .ALUT(n3197), .C0(address[1]), .Z(n3202));
    PFUMX i1263 (.BLUT(n3198), .ALUT(n3199), .C0(address[1]), .Z(n3203));
    PFUMX i1125 (.BLUT(n3057), .ALUT(n3058), .C0(address[1]), .Z(n3065));
    PFUMX i1126 (.BLUT(n3059), .ALUT(n3060), .C0(address[1]), .Z(n3066));
    PFUMX i1127 (.BLUT(n3061), .ALUT(n3062), .C0(address[1]), .Z(n3067));
    PFUMX i1128 (.BLUT(n3063), .ALUT(n3064), .C0(address[1]), .Z(n3068));
    PFUMX i1140 (.BLUT(n3072), .ALUT(n3073), .C0(address[1]), .Z(n3080));
    PFUMX i990 (.BLUT(n2922), .ALUT(n2923), .C0(address[1]), .Z(n2930));
    PFUMX i991 (.BLUT(n2924), .ALUT(n2925), .C0(address[1]), .Z(n2931));
    LUT4 \BUFF_5[[12__bdd_3_lut_1957  (.A(\BUFF[5] [12]), .B(\BUFF[7] [12]), 
         .C(address[1]), .Z(n3765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_5[[12__bdd_3_lut_1957 .init = 16'hcaca;
    LUT4 i1092_3_lut (.A(\BUFF[10] [0]), .B(\BUFF[11] [0]), .C(address[0]), 
         .Z(n3032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1092_3_lut.init = 16'hcaca;
    MUX21 i1523 (.D0(n2994), .D1(n2995), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[7]));
    PFUMX i1141 (.BLUT(n3074), .ALUT(n3075), .C0(address[1]), .Z(n3081));
    LUT4 \BUFF_5[[12__bdd_3_lut  (.A(\BUFF[4] [12]), .B(\BUFF[6] [12]), 
         .C(address[1]), .Z(n3766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_5[[12__bdd_3_lut .init = 16'hcaca;
    LUT4 \BUFF_0[[12__bdd_3_lut_1960  (.A(\BUFF[3] [12]), .B(\BUFF[1] [12]), 
         .C(address[1]), .Z(n3768)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam \BUFF_0[[12__bdd_3_lut_1960 .init = 16'hacac;
    LUT4 \BUFF_0[[12__bdd_3_lut  (.A(\BUFF[0] [12]), .B(\BUFF[2] [12]), 
         .C(address[1]), .Z(n3769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_0[[12__bdd_3_lut .init = 16'hcaca;
    PFUMX i1142 (.BLUT(n3076), .ALUT(n3077), .C0(address[1]), .Z(n3082));
    PFUMX i1143 (.BLUT(n3078), .ALUT(n3079), .C0(address[1]), .Z(n3083));
    MUX21 i1517 (.D0(n3054), .D1(n3055), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[4]));
    MUX21 i154033_i1 (.D0(n3750), .D1(n3764), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[1]));
    MUX21 i1499 (.D0(n2934), .D1(n3778), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[11]));
    MUX21 i1496 (.D0(n3084), .D1(n3085), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[2]));
    MUX21 i1524 (.D0(n2979), .D1(n2980), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[8]));
    MUX21 i1525 (.D0(n2964), .D1(n2965), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[9]));
    LUT4 \BUFF_13[[11__bdd_3_lut_1965  (.A(\BUFF[13] [11]), .B(\BUFF[15] [11]), 
         .C(address[1]), .Z(n3772)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_13[[11__bdd_3_lut_1965 .init = 16'hcaca;
    MUX21 i1518 (.D0(n3039), .D1(n3040), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[0]));
    LUT4 \BUFF_0[[1__bdd_3_lut  (.A(\BUFF[0] [1]), .B(\BUFF[2] [1]), .C(address[1]), 
         .Z(n3748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_0[[1__bdd_3_lut .init = 16'hcaca;
    MUX21 i1519 (.D0(n3189), .D1(n3190), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[14]));
    VHI i1973 (.Z(VCC_net));
    LUT4 \BUFF_13[[11__bdd_3_lut  (.A(\BUFF[12] [11]), .B(\BUFF[14] [11]), 
         .C(address[1]), .Z(n3773)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_13[[11__bdd_3_lut .init = 16'hcaca;
    MUX21 i1520 (.D0(n3024), .D1(n3025), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[5]));
    VLO i92 (.Z(GND_net));
    LUT4 \BUFF_5[[1__bdd_3_lut  (.A(\BUFF[4] [1]), .B(\BUFF[6] [1]), .C(address[1]), 
         .Z(n3745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_5[[1__bdd_3_lut .init = 16'hcaca;
    FD1P3AX BUFF_14__i0_i2 (.D(cpu_fpga_bus_d_out_2), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [2]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i2.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i3 (.D(cpu_fpga_bus_d_out_3), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [3]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i3.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i4 (.D(cpu_fpga_bus_d_out_4), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [4]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i4.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i5 (.D(cpu_fpga_bus_d_out_5), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [5]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i5.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i6 (.D(cpu_fpga_bus_d_out_6), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [6]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i6.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i7 (.D(cpu_fpga_bus_d_out_7), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [7]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i7.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i8 (.D(cpu_fpga_bus_d_out_8), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [8]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i8.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i9 (.D(cpu_fpga_bus_d_out_9), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [9]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i9.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i10 (.D(cpu_fpga_bus_d_out_10), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [10]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i10.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i11 (.D(cpu_fpga_bus_d_out_11), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [11]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i11.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i12 (.D(cpu_fpga_bus_d_out_12), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [12]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i12.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i13 (.D(cpu_fpga_bus_d_out_13), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [13]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i13.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i14 (.D(cpu_fpga_bus_d_out_14), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [14]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i14.GSR = "ENABLED";
    FD1P3AX BUFF_14__i0_i15 (.D(cpu_fpga_bus_d_out_15), .SP(cpu_fpga_clk_c_enable_260), 
            .CK(cpu_fpga_clk_c), .Q(\BUFF[14] [15]));   // /home/damiano/Documenti/Esami/Tesi/PUF/FPGA/impl1/source/top_level.vhd(37[3] 88[10])
    defparam BUFF_14__i0_i15.GSR = "ENABLED";
    LUT4 \BUFF_5[[1__bdd_3_lut_1933  (.A(\BUFF[5] [1]), .B(\BUFF[7] [1]), 
         .C(address[1]), .Z(n3744)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_5[[1__bdd_3_lut_1933 .init = 16'hcaca;
    MUX21 i153430_i1 (.D0(n3771), .D1(n3757), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[12]));
    L6MUX21 i1326 (.D0(n3264), .D1(n3265), .SD(\BUFF[0] [3]), .Z(fpga_io_gp_7__N_18[3]));
    LUT4 \BUFF_8[[11__bdd_3_lut_1968  (.A(\BUFF[11] [11]), .B(\BUFF[9] [11]), 
         .C(address[1]), .Z(n3775)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam \BUFF_8[[11__bdd_3_lut_1968 .init = 16'hacac;
    LUT4 \BUFF_8[[11__bdd_3_lut  (.A(\BUFF[8] [11]), .B(\BUFF[10] [11]), 
         .C(address[1]), .Z(n3776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \BUFF_8[[11__bdd_3_lut .init = 16'hcaca;
    LUT4 i1169_3_lut (.A(\BUFF[14] [0]), .B(\BUFF[15] [0]), .C(\BUFF[0] [0]), 
         .Z(n3109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1169_3_lut.init = 16'hcaca;
    MUX21 i1522 (.D0(n3009), .D1(n3010), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[6]));
    TSALL TSALL_INST (.TSALL(GND_net));
    L6MUX21 i1311 (.D0(n3249), .D1(n3250), .SD(\BUFF[0] [3]), .Z(fpga_io_gp_7__N_18[4]));
    LUT4 i1168_3_lut (.A(\BUFF[12] [0]), .B(\BUFF[13] [0]), .C(\BUFF[0] [0]), 
         .Z(n3108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1168_3_lut.init = 16'hcaca;
    LUT4 i1183_3_lut (.A(\BUFF[12] [6]), .B(\BUFF[13] [6]), .C(\BUFF[0] [0]), 
         .Z(n3123)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1183_3_lut.init = 16'hcaca;
    MUX21 i1515 (.D0(n3069), .D1(n3070), .SD(address[3]), .Z(cpu_fpga_bus_d_15__N_570[3]));
    L6MUX21 i1221 (.D0(n3159), .D1(n3160), .SD(\BUFF[0] [3]), .Z(fpga_io_gp_7__N_18[1]));
    LUT4 i1182_3_lut (.A(\BUFF[10] [6]), .B(\BUFF[11] [6]), .C(\BUFF[0] [0]), 
         .Z(n3122)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1182_3_lut.init = 16'hcaca;
    L6MUX21 i1296 (.D0(n3234), .D1(n3235), .SD(\BUFF[0] [3]), .Z(fpga_io_gp_7__N_18[7]));
    L6MUX21 i1206 (.D0(n3144), .D1(n3145), .SD(\BUFF[0] [3]), .Z(fpga_io_gp_7__N_18[5]));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    L6MUX21 i1191 (.D0(n3129), .D1(n3130), .SD(\BUFF[0] [3]), .Z(fpga_io_gp_7__N_18[6]));
    L6MUX21 i981 (.D0(n2919), .D1(n2920), .SD(\BUFF[0] [3]), .Z(fpga_io_gp_7__N_18[2]));
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

